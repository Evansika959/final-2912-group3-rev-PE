module 8b_mult (
    inout wire vss,
    inout wire vdd,
    inout wire a0_not,
    inout wire a0,
    inout wire a1_not,
    inout wire a1,
    inout wire a2_not,
    inout wire a2,
    inout wire a3_not,
    inout wire a3,
    inout wire a4_not,
    inout wire a4,
    inout wire a5_not,
    inout wire a5,
    inout wire a6_not,
    inout wire a6,
    inout wire a7_not,
    inout wire a7,
    inout wire b0_not,
    inout wire b0,
    inout wire b1_not,
    inout wire b1,
    inout wire p0,
    inout wire p0_not,
    inout wire p1,
    inout wire p1_not,
    inout wire b0_r1_b,
    inout wire b0_r1_b_not,
    inout wire b0_q0,
    inout wire b0_q0_not,
    inout wire b0_p0,
    inout wire b0_p0_not,
    inout wire b0_q1,
    inout wire b0_q1_not,
    inout wire b0_p1,
    inout wire b0_p1_not,
    inout wire b0_q2,
    inout wire b0_q2_not,
    inout wire b0_p2,
    inout wire b0_p2_not,
    inout wire b0_q3,
    inout wire b0_q3_not,
    inout wire b0_p3,
    inout wire b0_p3_not,
    inout wire b0_q4,
    inout wire b0_q4_not,
    inout wire b0_p4,
    inout wire b0_p4_not,
    inout wire b0_q5,
    inout wire b0_q5_not,
    inout wire b0_p5,
    inout wire b0_p5_not,
    inout wire b0_q6,
    inout wire b0_q6_not,
    inout wire b0_p6,
    inout wire b0_p6_not,
    inout wire b0_q7,
    inout wire b0_q7_not,
    inout wire b0_p7,
    inout wire b0_p7_not,
    inout wire b1_q7,
    inout wire b1_q7_not,
    inout wire b1_p7,
    inout wire b1_p7_not,
    inout wire b1_q6,
    inout wire b1_q6_not,
    inout wire b1_p6,
    inout wire b1_p6_not,
    inout wire b1_q5,
    inout wire b1_q5_not,
    inout wire b1_p5,
    inout wire b1_p5_not,
    inout wire b1_q4,
    inout wire b1_q4_not,
    inout wire b1_p4,
    inout wire b1_p4_not,
    inout wire b1_q3,
    inout wire b1_q3_not,
    inout wire b1_p3,
    inout wire b1_p3_not,
    inout wire b1_q2,
    inout wire b1_q2_not,
    inout wire b1_p2,
    inout wire b1_p2_not,
    inout wire b1_q1,
    inout wire b1_q1_not,
    inout wire b1_p1,
    inout wire b1_p1_not,
    inout wire b1_q0,
    inout wire b1_q0_not,
    inout wire b1_p0,
    inout wire b1_p0_not,
    inout wire b1_c0,
    inout wire b1_c0_not,
    inout wire b1_c1,
    inout wire b1_c1_not,
    inout wire b1_c2,
    inout wire b1_c2_not,
    inout wire b1_c3,
    inout wire b1_c3_not,
    inout wire b1_c4,
    inout wire b1_c4_not,
    inout wire b1_c5,
    inout wire b1_c5_not,
    inout wire b1_c6,
    inout wire b1_c6_not,
    inout wire b1_c7,
    inout wire b1_c7_not,
    inout wire b0_c7,
    inout wire b0_c7_not,
    inout wire b0_c6,
    inout wire b0_c6_not,
    inout wire b0_c5,
    inout wire b0_c5_not,
    inout wire b0_c4,
    inout wire b0_c4_not,
    inout wire b0_c3,
    inout wire b0_c3_not,
    inout wire b0_c2,
    inout wire b0_c2_not,
    inout wire b0_c1,
    inout wire b0_c1_not,
    inout wire b0_c0,
    inout wire b0_c0_not,
    inout wire b2_c0,
    inout wire b2_c0_not,
    inout wire b2_q0,
    inout wire b2_q0_not,
    inout wire b2_p0,
    inout wire b2_p0_not,
    inout wire b2_q1,
    inout wire b2_q1_not,
    inout wire b2_p1,
    inout wire b2_p1_not,
    inout wire b2_c1,
    inout wire b2_c1_not,
    inout wire b2_q2,
    inout wire b2_q2_not,
    inout wire b2_p2,
    inout wire b2_p2_not,
    inout wire b2_q3,
    inout wire b2_q3_not,
    inout wire b2_p3,
    inout wire b2_p3_not,
    inout wire b2_q4,
    inout wire b2_q4_not,
    inout wire b2_p4,
    inout wire b2_p4_not,
    inout wire b2_q5,
    inout wire b2_q5_not,
    inout wire b2_p5,
    inout wire b2_p5_not,
    inout wire b2_q6,
    inout wire b2_q6_not,
    inout wire b2_p6,
    inout wire b2_p6_not,
    inout wire b2_q7,
    inout wire b2_q7_not,
    inout wire b2_p7,
    inout wire b2_p7_not,
    inout wire b2_c3,
    inout wire b2_c3_not,
    inout wire b2_c4,
    inout wire b2_c4_not,
    inout wire b2_c5,
    inout wire b2_c5_not,
    inout wire b2_c6,
    inout wire b2_c6_not,
    inout wire b2_c7,
    inout wire b2_c7_not,
    inout wire x0_c0_f,
    inout wire x0_c0_f_not,
    inout wire x1_c0_f,
    inout wire x1_c0_f_not,
    inout wire x0_b0_f,
    inout wire x0_b0_f_not,
    inout wire x0_c0_b,
    inout wire x0_c0_b_not,
    inout wire b0_r2_b,
    inout wire b0_r2_b_not,
    inout wire b0_r3_b,
    inout wire b0_r3_b_not,
    inout wire b0_r4_b,
    inout wire b0_r4_b_not,
    inout wire b0_r5_b,
    inout wire b0_r5_b_not,
    inout wire b0_r6_b,
    inout wire b0_r6_b_not,
    inout wire b0_r7_b,
    inout wire b0_r7_b_not,
    inout wire x0_a7_f,
    inout wire x0_a7_f_not,
    inout wire x0_a7_b,
    inout wire x0_a7_b_not,
    inout wire x1_b0_f,
    inout wire x1_b0_f_not,
    inout wire p2,
    inout wire p2_not,
    inout wire x1_c0_b,
    inout wire x1_c0_b_not,
    inout wire b2_r0_b,
    inout wire b2_r0_b_not,
    inout wire b2_r1_b,
    inout wire b2_r1_b_not,
    inout wire b2_r2_b,
    inout wire b2_r2_b_not,
    inout wire b2_r3_b,
    inout wire b2_r3_b_not,
    inout wire b2_r4_b,
    inout wire b2_r4_b_not,
    inout wire b2_r5_b,
    inout wire b2_r5_b_not,
    inout wire b2_r6_b,
    inout wire b2_r6_b_not,
    inout wire b2_r7_b,
    inout wire b2_r7_b_not,
    inout wire b3_c0,
    inout wire b3_c0_not,
    inout wire b3_q0,
    inout wire b3_q0_not,
    inout wire b3_p0,
    inout wire b3_p0_not,
    inout wire b3_q1,
    inout wire b3_q1_not,
    inout wire b3_p1,
    inout wire b3_p1_not,
    inout wire b3_c1,
    inout wire b3_c1_not,
    inout wire b3_q2,
    inout wire b3_q2_not,
    inout wire b3_p2,
    inout wire b3_p2_not,
    inout wire b3_q3,
    inout wire b3_q3_not,
    inout wire b3_p3,
    inout wire b3_p3_not,
    inout wire b3_q4,
    inout wire b3_q4_not,
    inout wire b3_p4,
    inout wire b3_p4_not,
    inout wire b3_q5,
    inout wire b3_q5_not,
    inout wire b3_p5,
    inout wire b3_p5_not,
    inout wire b3_q6,
    inout wire b3_q6_not,
    inout wire b3_p6,
    inout wire b3_p6_not,
    inout wire b3_q7,
    inout wire b3_q7_not,
    inout wire b3_p7,
    inout wire b3_p7_not,
    inout wire b3_c3,
    inout wire b3_c3_not,
    inout wire b3_c4,
    inout wire b3_c4_not,
    inout wire b3_c5,
    inout wire b3_c5_not,
    inout wire b3_c6,
    inout wire b3_c6_not,
    inout wire b3_c7,
    inout wire b3_c7_not,
    inout wire x2_c0_f,
    inout wire x2_c0_f_not,
    inout wire x2_b0_f,
    inout wire x2_b0_f_not,
    inout wire p3,
    inout wire p3_not,
    inout wire x2_c0_b,
    inout wire x2_c0_b_not,
    inout wire b3_r0_b,
    inout wire b3_r0_b_not,
    inout wire b3_r1_b,
    inout wire b3_r1_b_not,
    inout wire b3_r2_b,
    inout wire b3_r2_b_not,
    inout wire b3_r3_b,
    inout wire b3_r3_b_not,
    inout wire b3_r4_b,
    inout wire b3_r4_b_not,
    inout wire b3_r5_b,
    inout wire b3_r5_b_not,
    inout wire b3_r6_b,
    inout wire b3_r6_b_not,
    inout wire b3_r7_b,
    inout wire b3_r7_b_not,
    inout wire b4_c0,
    inout wire b4_c0_not,
    inout wire b4_q0,
    inout wire b4_q0_not,
    inout wire b4_p0,
    inout wire b4_p0_not,
    inout wire b4_q1,
    inout wire b4_q1_not,
    inout wire b4_p1,
    inout wire b4_p1_not,
    inout wire b4_c1,
    inout wire b4_c1_not,
    inout wire b4_q2,
    inout wire b4_q2_not,
    inout wire b4_p2,
    inout wire b4_p2_not,
    inout wire b4_q3,
    inout wire b4_q3_not,
    inout wire b4_p3,
    inout wire b4_p3_not,
    inout wire b4_q4,
    inout wire b4_q4_not,
    inout wire b4_p4,
    inout wire b4_p4_not,
    inout wire b4_q5,
    inout wire b4_q5_not,
    inout wire b4_p5,
    inout wire b4_p5_not,
    inout wire b4_q6,
    inout wire b4_q6_not,
    inout wire b4_p6,
    inout wire b4_p6_not,
    inout wire b4_q7,
    inout wire b4_q7_not,
    inout wire b4_p7,
    inout wire b4_p7_not,
    inout wire b4_c3,
    inout wire b4_c3_not,
    inout wire b4_c4,
    inout wire b4_c4_not,
    inout wire b4_c5,
    inout wire b4_c5_not,
    inout wire b4_c6,
    inout wire b4_c6_not,
    inout wire b4_c7,
    inout wire b4_c7_not,
    inout wire x3_c0_f,
    inout wire x3_c0_f_not,
    inout wire x3_b0_f,
    inout wire x3_b0_f_not,
    inout wire p4,
    inout wire p4_not,
    inout wire x3_c0_b,
    inout wire x3_c0_b_not,
    inout wire b4_r0_b,
    inout wire b4_r0_b_not,
    inout wire b4_r1_b,
    inout wire b4_r1_b_not,
    inout wire b4_r2_b,
    inout wire b4_r2_b_not,
    inout wire b4_r3_b,
    inout wire b4_r3_b_not,
    inout wire b4_r4_b,
    inout wire b4_r4_b_not,
    inout wire b4_r5_b,
    inout wire b4_r5_b_not,
    inout wire b4_r6_b,
    inout wire b4_r6_b_not,
    inout wire b4_r7_b,
    inout wire b4_r7_b_not,
    inout wire b5_c0,
    inout wire b5_c0_not,
    inout wire b5_q0,
    inout wire b5_q0_not,
    inout wire b5_p0,
    inout wire b5_p0_not,
    inout wire b5_q1,
    inout wire b5_q1_not,
    inout wire b5_p1,
    inout wire b5_p1_not,
    inout wire b5_c1,
    inout wire b5_c1_not,
    inout wire b5_q2,
    inout wire b5_q2_not,
    inout wire b5_p2,
    inout wire b5_p2_not,
    inout wire b5_q3,
    inout wire b5_q3_not,
    inout wire b5_p3,
    inout wire b5_p3_not,
    inout wire b5_q4,
    inout wire b5_q4_not,
    inout wire b5_p4,
    inout wire b5_p4_not,
    inout wire b5_q5,
    inout wire b5_q5_not,
    inout wire b5_p5,
    inout wire b5_p5_not,
    inout wire b5_q6,
    inout wire b5_q6_not,
    inout wire b5_p6,
    inout wire b5_p6_not,
    inout wire b5_q7,
    inout wire b5_q7_not,
    inout wire b5_p7,
    inout wire b5_p7_not,
    inout wire b5_c3,
    inout wire b5_c3_not,
    inout wire b5_c4,
    inout wire b5_c4_not,
    inout wire b5_c5,
    inout wire b5_c5_not,
    inout wire b5_c6,
    inout wire b5_c6_not,
    inout wire b5_c7,
    inout wire b5_c7_not,
    inout wire x4_c0_f,
    inout wire x4_c0_f_not,
    inout wire x4_b0_f,
    inout wire x4_b0_f_not,
    inout wire p5,
    inout wire p5_not,
    inout wire x4_c0_b,
    inout wire x4_c0_b_not,
    inout wire b5_r0_b,
    inout wire b5_r0_b_not,
    inout wire b5_r1_b,
    inout wire b5_r1_b_not,
    inout wire b5_r2_b,
    inout wire b5_r2_b_not,
    inout wire b5_r3_b,
    inout wire b5_r3_b_not,
    inout wire b5_r4_b,
    inout wire b5_r4_b_not,
    inout wire b5_r5_b,
    inout wire b5_r5_b_not,
    inout wire b5_r6_b,
    inout wire b5_r6_b_not,
    inout wire b5_r7_b,
    inout wire b5_r7_b_not,
    inout wire b6_c0,
    inout wire b6_c0_not,
    inout wire b6_q0,
    inout wire b6_q0_not,
    inout wire b6_p0,
    inout wire b6_p0_not,
    inout wire b6_q1,
    inout wire b6_q1_not,
    inout wire b6_p1,
    inout wire b6_p1_not,
    inout wire b6_c1,
    inout wire b6_c1_not,
    inout wire b6_q2,
    inout wire b6_q2_not,
    inout wire b6_p2,
    inout wire b6_p2_not,
    inout wire b6_q3,
    inout wire b6_q3_not,
    inout wire b6_p3,
    inout wire b6_p3_not,
    inout wire b6_q4,
    inout wire b6_q4_not,
    inout wire b6_p4,
    inout wire b6_p4_not,
    inout wire b6_q5,
    inout wire b6_q5_not,
    inout wire b6_p5,
    inout wire b6_p5_not,
    inout wire b6_q6,
    inout wire b6_q6_not,
    inout wire b6_p6,
    inout wire b6_p6_not,
    inout wire b6_q7,
    inout wire b6_q7_not,
    inout wire b6_p7,
    inout wire b6_p7_not,
    inout wire b6_c3,
    inout wire b6_c3_not,
    inout wire b6_c4,
    inout wire b6_c4_not,
    inout wire b6_c5,
    inout wire b6_c5_not,
    inout wire b6_c6,
    inout wire b6_c6_not,
    inout wire b6_c7,
    inout wire b6_c7_not,
    inout wire x5_c0_f,
    inout wire x5_c0_f_not,
    inout wire x5_b0_f,
    inout wire x5_b0_f_not,
    inout wire p6,
    inout wire p6_not,
    inout wire x5_c0_b,
    inout wire x5_c0_b_not,
    inout wire b6_r0_b,
    inout wire b6_r0_b_not,
    inout wire b6_r1_b,
    inout wire b6_r1_b_not,
    inout wire b6_r2_b,
    inout wire b6_r2_b_not,
    inout wire b6_r3_b,
    inout wire b6_r3_b_not,
    inout wire b6_r4_b,
    inout wire b6_r4_b_not,
    inout wire b6_r5_b,
    inout wire b6_r5_b_not,
    inout wire b6_r6_b,
    inout wire b6_r6_b_not,
    inout wire b6_r7_b,
    inout wire b6_r7_b_not,
    inout wire b7_c0,
    inout wire b7_c0_not,
    inout wire b7_q0,
    inout wire b7_q0_not,
    inout wire b7_p0,
    inout wire b7_p0_not,
    inout wire b7_q1,
    inout wire b7_q1_not,
    inout wire b7_p1,
    inout wire b7_p1_not,
    inout wire b7_c1,
    inout wire b7_c1_not,
    inout wire b7_q2,
    inout wire b7_q2_not,
    inout wire b7_p2,
    inout wire b7_p2_not,
    inout wire b7_q3,
    inout wire b7_q3_not,
    inout wire b7_p3,
    inout wire b7_p3_not,
    inout wire b7_q4,
    inout wire b7_q4_not,
    inout wire b7_p4,
    inout wire b7_p4_not,
    inout wire b7_q5,
    inout wire b7_q5_not,
    inout wire b7_p5,
    inout wire b7_p5_not,
    inout wire b7_q6,
    inout wire b7_q6_not,
    inout wire b7_p6,
    inout wire b7_p6_not,
    inout wire b7_q7,
    inout wire b7_q7_not,
    inout wire b7_p7,
    inout wire b7_p7_not,
    inout wire b7_c3,
    inout wire b7_c3_not,
    inout wire b7_c4,
    inout wire b7_c4_not,
    inout wire b7_c5,
    inout wire b7_c5_not,
    inout wire b7_c6,
    inout wire b7_c6_not,
    inout wire b7_c7,
    inout wire b7_c7_not,
    inout wire x6_c0_f,
    inout wire x6_c0_f_not,
    inout wire x6_b0_f,
    inout wire x6_b0_f_not,
    inout wire p7,
    inout wire p7_not,
    inout wire x6_c0_b,
    inout wire x6_c0_b_not,
    inout wire b7_r0_b,
    inout wire b7_r0_b_not,
    inout wire b7_r1_b,
    inout wire b7_r1_b_not,
    inout wire b7_r2_b,
    inout wire b7_r2_b_not,
    inout wire b7_r3_b,
    inout wire b7_r3_b_not,
    inout wire b7_r4_b,
    inout wire b7_r4_b_not,
    inout wire b7_r5_b,
    inout wire b7_r5_b_not,
    inout wire b7_r6_b,
    inout wire b7_r6_b_not,
    inout wire b7_r7_b,
    inout wire b7_r7_b_not,
    inout wire p8,
    inout wire p8_not,
    inout wire p9,
    inout wire p9_not,
    inout wire p10,
    inout wire p10_not,
    inout wire p11,
    inout wire p11_not,
    inout wire p12,
    inout wire p12_not,
    inout wire p13,
    inout wire p13_not,
    inout wire p14,
    inout wire p14_not,
    inout wire p15,
    inout wire p15_not,
    inout wire b6_c2,
    inout wire b6_c2_not,
    inout wire b7_c2,
    inout wire b7_c2_not,
    inout wire b4_c2,
    inout wire b4_c2_not,
    inout wire b3_c2,
    inout wire b3_c2_not,
    inout wire b2_c2,
    inout wire b2_c2_not,
    inout wire b5_c2,
    inout wire b5_c2_not,
    inout wire b2_not,
    inout wire b2,
    inout wire b3_not,
    inout wire b3,
    inout wire b4_not,
    inout wire b4,
    inout wire b5_not,
    inout wire b5,
    inout wire b6_not,
    inout wire b6,
    inout wire b7_not,
    inout wire b7
);

endmodule