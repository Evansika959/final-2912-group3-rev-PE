(* blackbox *)
module fa_16b (
    inout wire VSS,
    inout wire VDD,
    inout wire z,
    inout wire z_not,
    inout wire c0_b,
    inout wire c0_not_b,
    inout wire c15_not,
    inout wire c15,
    inout wire s5_not,
    inout wire s5,
    inout wire s0_not,
    inout wire s0,
    inout wire s6_not,
    inout wire s6,
    inout wire s1_not,
    inout wire s1,
    inout wire s7_not,
    inout wire s7,
    inout wire s2_not,
    inout wire s2,
    inout wire s8_not,
    inout wire s8,
    inout wire s3_not,
    inout wire s3,
    inout wire s9_not,
    inout wire s9,
    inout wire s4_not,
    inout wire s4,
    inout wire s10_not,
    inout wire s10,
    inout wire s11_not,
    inout wire s11,
    inout wire s12_not,
    inout wire s12,
    inout wire s13_not,
    inout wire s13,
    inout wire s14_not,
    inout wire s14,
    inout wire s15_not,
    inout wire s15,
    inout wire c0_f,
    inout wire c0_f_not,
    inout wire a0_f,
    inout wire a0_not_f,
    inout wire b0,
    inout wire b0_not,
    inout wire a1_f,
    inout wire a1_not_f,
    inout wire b1,
    inout wire b1_not,
    inout wire a2_f,
    inout wire a2_not_f,
    inout wire b2,
    inout wire b2_not,
    inout wire a3_f,
    inout wire a3_not_f,
    inout wire b3,
    inout wire b3_not,
    inout wire a4_f,
    inout wire a4_not_f,
    inout wire b4,
    inout wire b4_not,
    inout wire a5_f,
    inout wire a5_not_f,
    inout wire b5,
    inout wire b5_not,
    inout wire a6_f,
    inout wire a6_not_f,
    inout wire b6,
    inout wire b6_not,
    inout wire a7_f,
    inout wire a7_not_f,
    inout wire b7,
    inout wire b7_not,
    inout wire a8_f,
    inout wire a8_not_f,
    inout wire b8,
    inout wire b8_not,
    inout wire a9_f,
    inout wire a9_not_f,
    inout wire b9,
    inout wire b9_not,
    inout wire a10_f,
    inout wire a10_not_f,
    inout wire b10,
    inout wire b10_not,
    inout wire a11_f,
    inout wire a11_not_f,
    inout wire b11,
    inout wire b11_not,
    inout wire a12_f,
    inout wire a12_not_f,
    inout wire b12,
    inout wire b12_not,
    inout wire a13_f,
    inout wire a13_not_f,
    inout wire b13,
    inout wire b13_not,
    inout wire a14_f,
    inout wire a14_not_f,
    inout wire b14,
    inout wire b14_not,
    inout wire a15_f,
    inout wire a15_not_f,
    inout wire b15,
    inout wire b15_not,
    inout wire a0_b,
    inout wire a0_not_b,
    inout wire a1_b,
    inout wire a1_not_b,
    inout wire a2_b,
    inout wire a2_not_b,
    inout wire a3_b,
    inout wire a3_not_b,
    inout wire a4_b,
    inout wire a4_not_b,
    inout wire a5_b,
    inout wire a5_not_b,
    inout wire a6_b,
    inout wire a6_not_b,
    inout wire a7_b,
    inout wire a7_not_b,
    inout wire a8_b,
    inout wire a8_not_b,
    inout wire a9_b,
    inout wire a9_not_b,
    inout wire a10_b,
    inout wire a10_not_b,
    inout wire a11_b,
    inout wire a11_not_b,
    inout wire a12_b,
    inout wire a12_not_b,
    inout wire a13_b,
    inout wire a13_not_b,
    inout wire a14_b,
    inout wire a14_not_b,
    inout wire a15_b,
    inout wire a15_not_b
);

endmodule